//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Formal Top-level netlist of Design: diffeq_paj_convert
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Dec  6 10:32:44 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module diffeq_paj_convert_top_formal_verification_random_tb;
// ----- Default clock port is added here since benchmark does not contain one -------
	reg [0:0] clk;

// ----- Shared inputs -------
	reg [0:0] Xinport_0_;
	reg [0:0] Xinport_1_;
	reg [0:0] Xinport_2_;
	reg [0:0] Xinport_3_;
	reg [0:0] Xinport_4_;
	reg [0:0] Xinport_5_;
	reg [0:0] Xinport_6_;
	reg [0:0] Xinport_7_;
	reg [0:0] Xinport_8_;
	reg [0:0] Xinport_9_;
	reg [0:0] Xinport_10_;
	reg [0:0] Xinport_11_;
	reg [0:0] Xinport_12_;
	reg [0:0] Xinport_13_;
	reg [0:0] Xinport_14_;
	reg [0:0] Xinport_15_;
	reg [0:0] Xinport_16_;
	reg [0:0] Xinport_17_;
	reg [0:0] Xinport_18_;
	reg [0:0] Xinport_19_;
	reg [0:0] Xinport_20_;
	reg [0:0] Xinport_21_;
	reg [0:0] Xinport_22_;
	reg [0:0] Xinport_23_;
	reg [0:0] Xinport_24_;
	reg [0:0] Xinport_25_;
	reg [0:0] Xinport_26_;
	reg [0:0] Xinport_27_;
	reg [0:0] Xinport_28_;
	reg [0:0] Xinport_29_;
	reg [0:0] Xinport_30_;
	reg [0:0] Xinport_31_;
	reg [0:0] Yinport_0_;
	reg [0:0] Yinport_1_;
	reg [0:0] Yinport_2_;
	reg [0:0] Yinport_3_;
	reg [0:0] Yinport_4_;
	reg [0:0] Yinport_5_;
	reg [0:0] Yinport_6_;
	reg [0:0] Yinport_7_;
	reg [0:0] Yinport_8_;
	reg [0:0] Yinport_9_;
	reg [0:0] Yinport_10_;
	reg [0:0] Yinport_11_;
	reg [0:0] Yinport_12_;
	reg [0:0] Yinport_13_;
	reg [0:0] Yinport_14_;
	reg [0:0] Yinport_15_;
	reg [0:0] Yinport_16_;
	reg [0:0] Yinport_17_;
	reg [0:0] Yinport_18_;
	reg [0:0] Yinport_19_;
	reg [0:0] Yinport_20_;
	reg [0:0] Yinport_21_;
	reg [0:0] Yinport_22_;
	reg [0:0] Yinport_23_;
	reg [0:0] Yinport_24_;
	reg [0:0] Yinport_25_;
	reg [0:0] Yinport_26_;
	reg [0:0] Yinport_27_;
	reg [0:0] Yinport_28_;
	reg [0:0] Yinport_29_;
	reg [0:0] Yinport_30_;
	reg [0:0] Yinport_31_;
	reg [0:0] Uinport_0_;
	reg [0:0] Uinport_1_;
	reg [0:0] Uinport_2_;
	reg [0:0] Uinport_3_;
	reg [0:0] Uinport_4_;
	reg [0:0] Uinport_5_;
	reg [0:0] Uinport_6_;
	reg [0:0] Uinport_7_;
	reg [0:0] Uinport_8_;
	reg [0:0] Uinport_9_;
	reg [0:0] Uinport_10_;
	reg [0:0] Uinport_11_;
	reg [0:0] Uinport_12_;
	reg [0:0] Uinport_13_;
	reg [0:0] Uinport_14_;
	reg [0:0] Uinport_15_;
	reg [0:0] Uinport_16_;
	reg [0:0] Uinport_17_;
	reg [0:0] Uinport_18_;
	reg [0:0] Uinport_19_;
	reg [0:0] Uinport_20_;
	reg [0:0] Uinport_21_;
	reg [0:0] Uinport_22_;
	reg [0:0] Uinport_23_;
	reg [0:0] Uinport_24_;
	reg [0:0] Uinport_25_;
	reg [0:0] Uinport_26_;
	reg [0:0] Uinport_27_;
	reg [0:0] Uinport_28_;
	reg [0:0] Uinport_29_;
	reg [0:0] Uinport_30_;
	reg [0:0] Uinport_31_;
	reg [0:0] Aport_0_;
	reg [0:0] Aport_1_;
	reg [0:0] Aport_2_;
	reg [0:0] Aport_3_;
	reg [0:0] Aport_4_;
	reg [0:0] Aport_5_;
	reg [0:0] Aport_6_;
	reg [0:0] Aport_7_;
	reg [0:0] Aport_8_;
	reg [0:0] Aport_9_;
	reg [0:0] Aport_10_;
	reg [0:0] Aport_11_;
	reg [0:0] Aport_12_;
	reg [0:0] Aport_13_;
	reg [0:0] Aport_14_;
	reg [0:0] Aport_15_;
	reg [0:0] Aport_16_;
	reg [0:0] Aport_17_;
	reg [0:0] Aport_18_;
	reg [0:0] Aport_19_;
	reg [0:0] Aport_20_;
	reg [0:0] Aport_21_;
	reg [0:0] Aport_22_;
	reg [0:0] Aport_23_;
	reg [0:0] Aport_24_;
	reg [0:0] Aport_25_;
	reg [0:0] Aport_26_;
	reg [0:0] Aport_27_;
	reg [0:0] Aport_28_;
	reg [0:0] Aport_29_;
	reg [0:0] Aport_30_;
	reg [0:0] Aport_31_;
	reg [0:0] DXport_0_;
	reg [0:0] DXport_1_;
	reg [0:0] DXport_2_;
	reg [0:0] DXport_3_;
	reg [0:0] DXport_4_;
	reg [0:0] DXport_5_;
	reg [0:0] DXport_6_;
	reg [0:0] DXport_7_;
	reg [0:0] DXport_8_;
	reg [0:0] DXport_9_;
	reg [0:0] DXport_10_;
	reg [0:0] DXport_11_;
	reg [0:0] DXport_12_;
	reg [0:0] DXport_13_;
	reg [0:0] DXport_14_;
	reg [0:0] DXport_15_;
	reg [0:0] DXport_16_;
	reg [0:0] DXport_17_;
	reg [0:0] DXport_18_;
	reg [0:0] DXport_19_;
	reg [0:0] DXport_20_;
	reg [0:0] DXport_21_;
	reg [0:0] DXport_22_;
	reg [0:0] DXport_23_;
	reg [0:0] DXport_24_;
	reg [0:0] DXport_25_;
	reg [0:0] DXport_26_;
	reg [0:0] DXport_27_;
	reg [0:0] DXport_28_;
	reg [0:0] DXport_29_;
	reg [0:0] DXport_30_;
	reg [0:0] DXport_31_;
	reg [0:0] reset;

// ----- FPGA fabric outputs -------
	wire [0:0] Xoutport_0__gfpga;
	wire [0:0] Xoutport_1__gfpga;
	wire [0:0] Xoutport_2__gfpga;
	wire [0:0] Xoutport_3__gfpga;
	wire [0:0] Xoutport_4__gfpga;
	wire [0:0] Xoutport_5__gfpga;
	wire [0:0] Xoutport_6__gfpga;
	wire [0:0] Xoutport_7__gfpga;
	wire [0:0] Xoutport_8__gfpga;
	wire [0:0] Xoutport_9__gfpga;
	wire [0:0] Xoutport_10__gfpga;
	wire [0:0] Xoutport_11__gfpga;
	wire [0:0] Xoutport_12__gfpga;
	wire [0:0] Xoutport_13__gfpga;
	wire [0:0] Xoutport_14__gfpga;
	wire [0:0] Xoutport_15__gfpga;
	wire [0:0] Xoutport_16__gfpga;
	wire [0:0] Xoutport_17__gfpga;
	wire [0:0] Xoutport_18__gfpga;
	wire [0:0] Xoutport_19__gfpga;
	wire [0:0] Xoutport_20__gfpga;
	wire [0:0] Xoutport_21__gfpga;
	wire [0:0] Xoutport_22__gfpga;
	wire [0:0] Xoutport_23__gfpga;
	wire [0:0] Xoutport_24__gfpga;
	wire [0:0] Xoutport_25__gfpga;
	wire [0:0] Xoutport_26__gfpga;
	wire [0:0] Xoutport_27__gfpga;
	wire [0:0] Xoutport_28__gfpga;
	wire [0:0] Xoutport_29__gfpga;
	wire [0:0] Xoutport_30__gfpga;
	wire [0:0] Xoutport_31__gfpga;
	wire [0:0] Youtport_0__gfpga;
	wire [0:0] Youtport_1__gfpga;
	wire [0:0] Youtport_2__gfpga;
	wire [0:0] Youtport_3__gfpga;
	wire [0:0] Youtport_4__gfpga;
	wire [0:0] Youtport_5__gfpga;
	wire [0:0] Youtport_6__gfpga;
	wire [0:0] Youtport_7__gfpga;
	wire [0:0] Youtport_8__gfpga;
	wire [0:0] Youtport_9__gfpga;
	wire [0:0] Youtport_10__gfpga;
	wire [0:0] Youtport_11__gfpga;
	wire [0:0] Youtport_12__gfpga;
	wire [0:0] Youtport_13__gfpga;
	wire [0:0] Youtport_14__gfpga;
	wire [0:0] Youtport_15__gfpga;
	wire [0:0] Youtport_16__gfpga;
	wire [0:0] Youtport_17__gfpga;
	wire [0:0] Youtport_18__gfpga;
	wire [0:0] Youtport_19__gfpga;
	wire [0:0] Youtport_20__gfpga;
	wire [0:0] Youtport_21__gfpga;
	wire [0:0] Youtport_22__gfpga;
	wire [0:0] Youtport_23__gfpga;
	wire [0:0] Youtport_24__gfpga;
	wire [0:0] Youtport_25__gfpga;
	wire [0:0] Youtport_26__gfpga;
	wire [0:0] Youtport_27__gfpga;
	wire [0:0] Youtport_28__gfpga;
	wire [0:0] Youtport_29__gfpga;
	wire [0:0] Youtport_30__gfpga;
	wire [0:0] Youtport_31__gfpga;
	wire [0:0] Uoutport_0__gfpga;
	wire [0:0] Uoutport_1__gfpga;
	wire [0:0] Uoutport_2__gfpga;
	wire [0:0] Uoutport_3__gfpga;
	wire [0:0] Uoutport_4__gfpga;
	wire [0:0] Uoutport_5__gfpga;
	wire [0:0] Uoutport_6__gfpga;
	wire [0:0] Uoutport_7__gfpga;
	wire [0:0] Uoutport_8__gfpga;
	wire [0:0] Uoutport_9__gfpga;
	wire [0:0] Uoutport_10__gfpga;
	wire [0:0] Uoutport_11__gfpga;
	wire [0:0] Uoutport_12__gfpga;
	wire [0:0] Uoutport_13__gfpga;
	wire [0:0] Uoutport_14__gfpga;
	wire [0:0] Uoutport_15__gfpga;
	wire [0:0] Uoutport_16__gfpga;
	wire [0:0] Uoutport_17__gfpga;
	wire [0:0] Uoutport_18__gfpga;
	wire [0:0] Uoutport_19__gfpga;
	wire [0:0] Uoutport_20__gfpga;
	wire [0:0] Uoutport_21__gfpga;
	wire [0:0] Uoutport_22__gfpga;
	wire [0:0] Uoutport_23__gfpga;
	wire [0:0] Uoutport_24__gfpga;
	wire [0:0] Uoutport_25__gfpga;
	wire [0:0] Uoutport_26__gfpga;
	wire [0:0] Uoutport_27__gfpga;
	wire [0:0] Uoutport_28__gfpga;
	wire [0:0] Uoutport_29__gfpga;
	wire [0:0] Uoutport_30__gfpga;
	wire [0:0] Uoutport_31__gfpga;

// ----- Benchmark outputs -------
	wire [0:0] Xoutport_0__bench;
	wire [0:0] Xoutport_1__bench;
	wire [0:0] Xoutport_2__bench;
	wire [0:0] Xoutport_3__bench;
	wire [0:0] Xoutport_4__bench;
	wire [0:0] Xoutport_5__bench;
	wire [0:0] Xoutport_6__bench;
	wire [0:0] Xoutport_7__bench;
	wire [0:0] Xoutport_8__bench;
	wire [0:0] Xoutport_9__bench;
	wire [0:0] Xoutport_10__bench;
	wire [0:0] Xoutport_11__bench;
	wire [0:0] Xoutport_12__bench;
	wire [0:0] Xoutport_13__bench;
	wire [0:0] Xoutport_14__bench;
	wire [0:0] Xoutport_15__bench;
	wire [0:0] Xoutport_16__bench;
	wire [0:0] Xoutport_17__bench;
	wire [0:0] Xoutport_18__bench;
	wire [0:0] Xoutport_19__bench;
	wire [0:0] Xoutport_20__bench;
	wire [0:0] Xoutport_21__bench;
	wire [0:0] Xoutport_22__bench;
	wire [0:0] Xoutport_23__bench;
	wire [0:0] Xoutport_24__bench;
	wire [0:0] Xoutport_25__bench;
	wire [0:0] Xoutport_26__bench;
	wire [0:0] Xoutport_27__bench;
	wire [0:0] Xoutport_28__bench;
	wire [0:0] Xoutport_29__bench;
	wire [0:0] Xoutport_30__bench;
	wire [0:0] Xoutport_31__bench;
	wire [0:0] Youtport_0__bench;
	wire [0:0] Youtport_1__bench;
	wire [0:0] Youtport_2__bench;
	wire [0:0] Youtport_3__bench;
	wire [0:0] Youtport_4__bench;
	wire [0:0] Youtport_5__bench;
	wire [0:0] Youtport_6__bench;
	wire [0:0] Youtport_7__bench;
	wire [0:0] Youtport_8__bench;
	wire [0:0] Youtport_9__bench;
	wire [0:0] Youtport_10__bench;
	wire [0:0] Youtport_11__bench;
	wire [0:0] Youtport_12__bench;
	wire [0:0] Youtport_13__bench;
	wire [0:0] Youtport_14__bench;
	wire [0:0] Youtport_15__bench;
	wire [0:0] Youtport_16__bench;
	wire [0:0] Youtport_17__bench;
	wire [0:0] Youtport_18__bench;
	wire [0:0] Youtport_19__bench;
	wire [0:0] Youtport_20__bench;
	wire [0:0] Youtport_21__bench;
	wire [0:0] Youtport_22__bench;
	wire [0:0] Youtport_23__bench;
	wire [0:0] Youtport_24__bench;
	wire [0:0] Youtport_25__bench;
	wire [0:0] Youtport_26__bench;
	wire [0:0] Youtport_27__bench;
	wire [0:0] Youtport_28__bench;
	wire [0:0] Youtport_29__bench;
	wire [0:0] Youtport_30__bench;
	wire [0:0] Youtport_31__bench;
	wire [0:0] Uoutport_0__bench;
	wire [0:0] Uoutport_1__bench;
	wire [0:0] Uoutport_2__bench;
	wire [0:0] Uoutport_3__bench;
	wire [0:0] Uoutport_4__bench;
	wire [0:0] Uoutport_5__bench;
	wire [0:0] Uoutport_6__bench;
	wire [0:0] Uoutport_7__bench;
	wire [0:0] Uoutport_8__bench;
	wire [0:0] Uoutport_9__bench;
	wire [0:0] Uoutport_10__bench;
	wire [0:0] Uoutport_11__bench;
	wire [0:0] Uoutport_12__bench;
	wire [0:0] Uoutport_13__bench;
	wire [0:0] Uoutport_14__bench;
	wire [0:0] Uoutport_15__bench;
	wire [0:0] Uoutport_16__bench;
	wire [0:0] Uoutport_17__bench;
	wire [0:0] Uoutport_18__bench;
	wire [0:0] Uoutport_19__bench;
	wire [0:0] Uoutport_20__bench;
	wire [0:0] Uoutport_21__bench;
	wire [0:0] Uoutport_22__bench;
	wire [0:0] Uoutport_23__bench;
	wire [0:0] Uoutport_24__bench;
	wire [0:0] Uoutport_25__bench;
	wire [0:0] Uoutport_26__bench;
	wire [0:0] Uoutport_27__bench;
	wire [0:0] Uoutport_28__bench;
	wire [0:0] Uoutport_29__bench;
	wire [0:0] Uoutport_30__bench;
	wire [0:0] Uoutport_31__bench;

// ----- Output vectors checking flags -------
	reg [0:0] Xoutport_0__flag;
	reg [0:0] Xoutport_1__flag;
	reg [0:0] Xoutport_2__flag;
	reg [0:0] Xoutport_3__flag;
	reg [0:0] Xoutport_4__flag;
	reg [0:0] Xoutport_5__flag;
	reg [0:0] Xoutport_6__flag;
	reg [0:0] Xoutport_7__flag;
	reg [0:0] Xoutport_8__flag;
	reg [0:0] Xoutport_9__flag;
	reg [0:0] Xoutport_10__flag;
	reg [0:0] Xoutport_11__flag;
	reg [0:0] Xoutport_12__flag;
	reg [0:0] Xoutport_13__flag;
	reg [0:0] Xoutport_14__flag;
	reg [0:0] Xoutport_15__flag;
	reg [0:0] Xoutport_16__flag;
	reg [0:0] Xoutport_17__flag;
	reg [0:0] Xoutport_18__flag;
	reg [0:0] Xoutport_19__flag;
	reg [0:0] Xoutport_20__flag;
	reg [0:0] Xoutport_21__flag;
	reg [0:0] Xoutport_22__flag;
	reg [0:0] Xoutport_23__flag;
	reg [0:0] Xoutport_24__flag;
	reg [0:0] Xoutport_25__flag;
	reg [0:0] Xoutport_26__flag;
	reg [0:0] Xoutport_27__flag;
	reg [0:0] Xoutport_28__flag;
	reg [0:0] Xoutport_29__flag;
	reg [0:0] Xoutport_30__flag;
	reg [0:0] Xoutport_31__flag;
	reg [0:0] Youtport_0__flag;
	reg [0:0] Youtport_1__flag;
	reg [0:0] Youtport_2__flag;
	reg [0:0] Youtport_3__flag;
	reg [0:0] Youtport_4__flag;
	reg [0:0] Youtport_5__flag;
	reg [0:0] Youtport_6__flag;
	reg [0:0] Youtport_7__flag;
	reg [0:0] Youtport_8__flag;
	reg [0:0] Youtport_9__flag;
	reg [0:0] Youtport_10__flag;
	reg [0:0] Youtport_11__flag;
	reg [0:0] Youtport_12__flag;
	reg [0:0] Youtport_13__flag;
	reg [0:0] Youtport_14__flag;
	reg [0:0] Youtport_15__flag;
	reg [0:0] Youtport_16__flag;
	reg [0:0] Youtport_17__flag;
	reg [0:0] Youtport_18__flag;
	reg [0:0] Youtport_19__flag;
	reg [0:0] Youtport_20__flag;
	reg [0:0] Youtport_21__flag;
	reg [0:0] Youtport_22__flag;
	reg [0:0] Youtport_23__flag;
	reg [0:0] Youtport_24__flag;
	reg [0:0] Youtport_25__flag;
	reg [0:0] Youtport_26__flag;
	reg [0:0] Youtport_27__flag;
	reg [0:0] Youtport_28__flag;
	reg [0:0] Youtport_29__flag;
	reg [0:0] Youtport_30__flag;
	reg [0:0] Youtport_31__flag;
	reg [0:0] Uoutport_0__flag;
	reg [0:0] Uoutport_1__flag;
	reg [0:0] Uoutport_2__flag;
	reg [0:0] Uoutport_3__flag;
	reg [0:0] Uoutport_4__flag;
	reg [0:0] Uoutport_5__flag;
	reg [0:0] Uoutport_6__flag;
	reg [0:0] Uoutport_7__flag;
	reg [0:0] Uoutport_8__flag;
	reg [0:0] Uoutport_9__flag;
	reg [0:0] Uoutport_10__flag;
	reg [0:0] Uoutport_11__flag;
	reg [0:0] Uoutport_12__flag;
	reg [0:0] Uoutport_13__flag;
	reg [0:0] Uoutport_14__flag;
	reg [0:0] Uoutport_15__flag;
	reg [0:0] Uoutport_16__flag;
	reg [0:0] Uoutport_17__flag;
	reg [0:0] Uoutport_18__flag;
	reg [0:0] Uoutport_19__flag;
	reg [0:0] Uoutport_20__flag;
	reg [0:0] Uoutport_21__flag;
	reg [0:0] Uoutport_22__flag;
	reg [0:0] Uoutport_23__flag;
	reg [0:0] Uoutport_24__flag;
	reg [0:0] Uoutport_25__flag;
	reg [0:0] Uoutport_26__flag;
	reg [0:0] Uoutport_27__flag;
	reg [0:0] Uoutport_28__flag;
	reg [0:0] Uoutport_29__flag;
	reg [0:0] Uoutport_30__flag;
	reg [0:0] Uoutport_31__flag;

// ----- Error counter -------
	integer nb_error= 0;

// ----- FPGA fabric instanciation -------
	diffeq_paj_convert_top_formal_verification FPGA_DUT(
		Xinport_0_,
		Xinport_1_,
		Xinport_2_,
		Xinport_3_,
		Xinport_4_,
		Xinport_5_,
		Xinport_6_,
		Xinport_7_,
		Xinport_8_,
		Xinport_9_,
		Xinport_10_,
		Xinport_11_,
		Xinport_12_,
		Xinport_13_,
		Xinport_14_,
		Xinport_15_,
		Xinport_16_,
		Xinport_17_,
		Xinport_18_,
		Xinport_19_,
		Xinport_20_,
		Xinport_21_,
		Xinport_22_,
		Xinport_23_,
		Xinport_24_,
		Xinport_25_,
		Xinport_26_,
		Xinport_27_,
		Xinport_28_,
		Xinport_29_,
		Xinport_30_,
		Xinport_31_,
		Yinport_0_,
		Yinport_1_,
		Yinport_2_,
		Yinport_3_,
		Yinport_4_,
		Yinport_5_,
		Yinport_6_,
		Yinport_7_,
		Yinport_8_,
		Yinport_9_,
		Yinport_10_,
		Yinport_11_,
		Yinport_12_,
		Yinport_13_,
		Yinport_14_,
		Yinport_15_,
		Yinport_16_,
		Yinport_17_,
		Yinport_18_,
		Yinport_19_,
		Yinport_20_,
		Yinport_21_,
		Yinport_22_,
		Yinport_23_,
		Yinport_24_,
		Yinport_25_,
		Yinport_26_,
		Yinport_27_,
		Yinport_28_,
		Yinport_29_,
		Yinport_30_,
		Yinport_31_,
		Uinport_0_,
		Uinport_1_,
		Uinport_2_,
		Uinport_3_,
		Uinport_4_,
		Uinport_5_,
		Uinport_6_,
		Uinport_7_,
		Uinport_8_,
		Uinport_9_,
		Uinport_10_,
		Uinport_11_,
		Uinport_12_,
		Uinport_13_,
		Uinport_14_,
		Uinport_15_,
		Uinport_16_,
		Uinport_17_,
		Uinport_18_,
		Uinport_19_,
		Uinport_20_,
		Uinport_21_,
		Uinport_22_,
		Uinport_23_,
		Uinport_24_,
		Uinport_25_,
		Uinport_26_,
		Uinport_27_,
		Uinport_28_,
		Uinport_29_,
		Uinport_30_,
		Uinport_31_,
		Aport_0_,
		Aport_1_,
		Aport_2_,
		Aport_3_,
		Aport_4_,
		Aport_5_,
		Aport_6_,
		Aport_7_,
		Aport_8_,
		Aport_9_,
		Aport_10_,
		Aport_11_,
		Aport_12_,
		Aport_13_,
		Aport_14_,
		Aport_15_,
		Aport_16_,
		Aport_17_,
		Aport_18_,
		Aport_19_,
		Aport_20_,
		Aport_21_,
		Aport_22_,
		Aport_23_,
		Aport_24_,
		Aport_25_,
		Aport_26_,
		Aport_27_,
		Aport_28_,
		Aport_29_,
		Aport_30_,
		Aport_31_,
		DXport_0_,
		DXport_1_,
		DXport_2_,
		DXport_3_,
		DXport_4_,
		DXport_5_,
		DXport_6_,
		DXport_7_,
		DXport_8_,
		DXport_9_,
		DXport_10_,
		DXport_11_,
		DXport_12_,
		DXport_13_,
		DXport_14_,
		DXport_15_,
		DXport_16_,
		DXport_17_,
		DXport_18_,
		DXport_19_,
		DXport_20_,
		DXport_21_,
		DXport_22_,
		DXport_23_,
		DXport_24_,
		DXport_25_,
		DXport_26_,
		DXport_27_,
		DXport_28_,
		DXport_29_,
		DXport_30_,
		DXport_31_,
		clk,
		reset,
		Xoutport_0__gfpga,
		Xoutport_1__gfpga,
		Xoutport_2__gfpga,
		Xoutport_3__gfpga,
		Xoutport_4__gfpga,
		Xoutport_5__gfpga,
		Xoutport_6__gfpga,
		Xoutport_7__gfpga,
		Xoutport_8__gfpga,
		Xoutport_9__gfpga,
		Xoutport_10__gfpga,
		Xoutport_11__gfpga,
		Xoutport_12__gfpga,
		Xoutport_13__gfpga,
		Xoutport_14__gfpga,
		Xoutport_15__gfpga,
		Xoutport_16__gfpga,
		Xoutport_17__gfpga,
		Xoutport_18__gfpga,
		Xoutport_19__gfpga,
		Xoutport_20__gfpga,
		Xoutport_21__gfpga,
		Xoutport_22__gfpga,
		Xoutport_23__gfpga,
		Xoutport_24__gfpga,
		Xoutport_25__gfpga,
		Xoutport_26__gfpga,
		Xoutport_27__gfpga,
		Xoutport_28__gfpga,
		Xoutport_29__gfpga,
		Xoutport_30__gfpga,
		Xoutport_31__gfpga,
		Youtport_0__gfpga,
		Youtport_1__gfpga,
		Youtport_2__gfpga,
		Youtport_3__gfpga,
		Youtport_4__gfpga,
		Youtport_5__gfpga,
		Youtport_6__gfpga,
		Youtport_7__gfpga,
		Youtport_8__gfpga,
		Youtport_9__gfpga,
		Youtport_10__gfpga,
		Youtport_11__gfpga,
		Youtport_12__gfpga,
		Youtport_13__gfpga,
		Youtport_14__gfpga,
		Youtport_15__gfpga,
		Youtport_16__gfpga,
		Youtport_17__gfpga,
		Youtport_18__gfpga,
		Youtport_19__gfpga,
		Youtport_20__gfpga,
		Youtport_21__gfpga,
		Youtport_22__gfpga,
		Youtport_23__gfpga,
		Youtport_24__gfpga,
		Youtport_25__gfpga,
		Youtport_26__gfpga,
		Youtport_27__gfpga,
		Youtport_28__gfpga,
		Youtport_29__gfpga,
		Youtport_30__gfpga,
		Youtport_31__gfpga,
		Uoutport_0__gfpga,
		Uoutport_1__gfpga,
		Uoutport_2__gfpga,
		Uoutport_3__gfpga,
		Uoutport_4__gfpga,
		Uoutport_5__gfpga,
		Uoutport_6__gfpga,
		Uoutport_7__gfpga,
		Uoutport_8__gfpga,
		Uoutport_9__gfpga,
		Uoutport_10__gfpga,
		Uoutport_11__gfpga,
		Uoutport_12__gfpga,
		Uoutport_13__gfpga,
		Uoutport_14__gfpga,
		Uoutport_15__gfpga,
		Uoutport_16__gfpga,
		Uoutport_17__gfpga,
		Uoutport_18__gfpga,
		Uoutport_19__gfpga,
		Uoutport_20__gfpga,
		Uoutport_21__gfpga,
		Uoutport_22__gfpga,
		Uoutport_23__gfpga,
		Uoutport_24__gfpga,
		Uoutport_25__gfpga,
		Uoutport_26__gfpga,
		Uoutport_27__gfpga,
		Uoutport_28__gfpga,
		Uoutport_29__gfpga,
		Uoutport_30__gfpga,
		Uoutport_31__gfpga
	);
// ----- End FPGA Fabric Instanication -------

// ----- Reference Benchmark Instanication -------
	diffeq_paj_convert REF_DUT(
		Xinport_0_,
		Xinport_1_,
		Xinport_2_,
		Xinport_3_,
		Xinport_4_,
		Xinport_5_,
		Xinport_6_,
		Xinport_7_,
		Xinport_8_,
		Xinport_9_,
		Xinport_10_,
		Xinport_11_,
		Xinport_12_,
		Xinport_13_,
		Xinport_14_,
		Xinport_15_,
		Xinport_16_,
		Xinport_17_,
		Xinport_18_,
		Xinport_19_,
		Xinport_20_,
		Xinport_21_,
		Xinport_22_,
		Xinport_23_,
		Xinport_24_,
		Xinport_25_,
		Xinport_26_,
		Xinport_27_,
		Xinport_28_,
		Xinport_29_,
		Xinport_30_,
		Xinport_31_,
		Yinport_0_,
		Yinport_1_,
		Yinport_2_,
		Yinport_3_,
		Yinport_4_,
		Yinport_5_,
		Yinport_6_,
		Yinport_7_,
		Yinport_8_,
		Yinport_9_,
		Yinport_10_,
		Yinport_11_,
		Yinport_12_,
		Yinport_13_,
		Yinport_14_,
		Yinport_15_,
		Yinport_16_,
		Yinport_17_,
		Yinport_18_,
		Yinport_19_,
		Yinport_20_,
		Yinport_21_,
		Yinport_22_,
		Yinport_23_,
		Yinport_24_,
		Yinport_25_,
		Yinport_26_,
		Yinport_27_,
		Yinport_28_,
		Yinport_29_,
		Yinport_30_,
		Yinport_31_,
		Uinport_0_,
		Uinport_1_,
		Uinport_2_,
		Uinport_3_,
		Uinport_4_,
		Uinport_5_,
		Uinport_6_,
		Uinport_7_,
		Uinport_8_,
		Uinport_9_,
		Uinport_10_,
		Uinport_11_,
		Uinport_12_,
		Uinport_13_,
		Uinport_14_,
		Uinport_15_,
		Uinport_16_,
		Uinport_17_,
		Uinport_18_,
		Uinport_19_,
		Uinport_20_,
		Uinport_21_,
		Uinport_22_,
		Uinport_23_,
		Uinport_24_,
		Uinport_25_,
		Uinport_26_,
		Uinport_27_,
		Uinport_28_,
		Uinport_29_,
		Uinport_30_,
		Uinport_31_,
		Aport_0_,
		Aport_1_,
		Aport_2_,
		Aport_3_,
		Aport_4_,
		Aport_5_,
		Aport_6_,
		Aport_7_,
		Aport_8_,
		Aport_9_,
		Aport_10_,
		Aport_11_,
		Aport_12_,
		Aport_13_,
		Aport_14_,
		Aport_15_,
		Aport_16_,
		Aport_17_,
		Aport_18_,
		Aport_19_,
		Aport_20_,
		Aport_21_,
		Aport_22_,
		Aport_23_,
		Aport_24_,
		Aport_25_,
		Aport_26_,
		Aport_27_,
		Aport_28_,
		Aport_29_,
		Aport_30_,
		Aport_31_,
		DXport_0_,
		DXport_1_,
		DXport_2_,
		DXport_3_,
		DXport_4_,
		DXport_5_,
		DXport_6_,
		DXport_7_,
		DXport_8_,
		DXport_9_,
		DXport_10_,
		DXport_11_,
		DXport_12_,
		DXport_13_,
		DXport_14_,
		DXport_15_,
		DXport_16_,
		DXport_17_,
		DXport_18_,
		DXport_19_,
		DXport_20_,
		DXport_21_,
		DXport_22_,
		DXport_23_,
		DXport_24_,
		DXport_25_,
		DXport_26_,
		DXport_27_,
		DXport_28_,
		DXport_29_,
		DXport_30_,
		DXport_31_,
		clk,
		reset,
		Xoutport_0__bench,
		Xoutport_1__bench,
		Xoutport_2__bench,
		Xoutport_3__bench,
		Xoutport_4__bench,
		Xoutport_5__bench,
		Xoutport_6__bench,
		Xoutport_7__bench,
		Xoutport_8__bench,
		Xoutport_9__bench,
		Xoutport_10__bench,
		Xoutport_11__bench,
		Xoutport_12__bench,
		Xoutport_13__bench,
		Xoutport_14__bench,
		Xoutport_15__bench,
		Xoutport_16__bench,
		Xoutport_17__bench,
		Xoutport_18__bench,
		Xoutport_19__bench,
		Xoutport_20__bench,
		Xoutport_21__bench,
		Xoutport_22__bench,
		Xoutport_23__bench,
		Xoutport_24__bench,
		Xoutport_25__bench,
		Xoutport_26__bench,
		Xoutport_27__bench,
		Xoutport_28__bench,
		Xoutport_29__bench,
		Xoutport_30__bench,
		Xoutport_31__bench,
		Youtport_0__bench,
		Youtport_1__bench,
		Youtport_2__bench,
		Youtport_3__bench,
		Youtport_4__bench,
		Youtport_5__bench,
		Youtport_6__bench,
		Youtport_7__bench,
		Youtport_8__bench,
		Youtport_9__bench,
		Youtport_10__bench,
		Youtport_11__bench,
		Youtport_12__bench,
		Youtport_13__bench,
		Youtport_14__bench,
		Youtport_15__bench,
		Youtport_16__bench,
		Youtport_17__bench,
		Youtport_18__bench,
		Youtport_19__bench,
		Youtport_20__bench,
		Youtport_21__bench,
		Youtport_22__bench,
		Youtport_23__bench,
		Youtport_24__bench,
		Youtport_25__bench,
		Youtport_26__bench,
		Youtport_27__bench,
		Youtport_28__bench,
		Youtport_29__bench,
		Youtport_30__bench,
		Youtport_31__bench,
		Uoutport_0__bench,
		Uoutport_1__bench,
		Uoutport_2__bench,
		Uoutport_3__bench,
		Uoutport_4__bench,
		Uoutport_5__bench,
		Uoutport_6__bench,
		Uoutport_7__bench,
		Uoutport_8__bench,
		Uoutport_9__bench,
		Uoutport_10__bench,
		Uoutport_11__bench,
		Uoutport_12__bench,
		Uoutport_13__bench,
		Uoutport_14__bench,
		Uoutport_15__bench,
		Uoutport_16__bench,
		Uoutport_17__bench,
		Uoutport_18__bench,
		Uoutport_19__bench,
		Uoutport_20__bench,
		Uoutport_21__bench,
		Uoutport_22__bench,
		Uoutport_23__bench,
		Uoutport_24__bench,
		Uoutport_25__bench,
		Uoutport_26__bench,
		Uoutport_27__bench,
		Uoutport_28__bench,
		Uoutport_29__bench,
		Uoutport_30__bench,
		Uoutport_31__bench
	);
// ----- End reference Benchmark Instanication -------

// ----- Clock 'clk' Initialization -------
	initial begin
		clk[0] <= 1'b0;
		while(1) begin
			#1
			clk[0] <= !clk[0];
		end
	end

// ----- Begin reset signal generation -----
// ----- End reset signal generation -----

// ----- Input Initialization -------
	initial begin
		Xinport_0_ <= 1'b0;
		Xinport_1_ <= 1'b0;
		Xinport_2_ <= 1'b0;
		Xinport_3_ <= 1'b0;
		Xinport_4_ <= 1'b0;
		Xinport_5_ <= 1'b0;
		Xinport_6_ <= 1'b0;
		Xinport_7_ <= 1'b0;
		Xinport_8_ <= 1'b0;
		Xinport_9_ <= 1'b0;
		Xinport_10_ <= 1'b0;
		Xinport_11_ <= 1'b0;
		Xinport_12_ <= 1'b0;
		Xinport_13_ <= 1'b0;
		Xinport_14_ <= 1'b0;
		Xinport_15_ <= 1'b0;
		Xinport_16_ <= 1'b0;
		Xinport_17_ <= 1'b0;
		Xinport_18_ <= 1'b0;
		Xinport_19_ <= 1'b0;
		Xinport_20_ <= 1'b0;
		Xinport_21_ <= 1'b0;
		Xinport_22_ <= 1'b0;
		Xinport_23_ <= 1'b0;
		Xinport_24_ <= 1'b0;
		Xinport_25_ <= 1'b0;
		Xinport_26_ <= 1'b0;
		Xinport_27_ <= 1'b0;
		Xinport_28_ <= 1'b0;
		Xinport_29_ <= 1'b0;
		Xinport_30_ <= 1'b0;
		Xinport_31_ <= 1'b0;
		Yinport_0_ <= 1'b0;
		Yinport_1_ <= 1'b0;
		Yinport_2_ <= 1'b0;
		Yinport_3_ <= 1'b0;
		Yinport_4_ <= 1'b0;
		Yinport_5_ <= 1'b0;
		Yinport_6_ <= 1'b0;
		Yinport_7_ <= 1'b0;
		Yinport_8_ <= 1'b0;
		Yinport_9_ <= 1'b0;
		Yinport_10_ <= 1'b0;
		Yinport_11_ <= 1'b0;
		Yinport_12_ <= 1'b0;
		Yinport_13_ <= 1'b0;
		Yinport_14_ <= 1'b0;
		Yinport_15_ <= 1'b0;
		Yinport_16_ <= 1'b0;
		Yinport_17_ <= 1'b0;
		Yinport_18_ <= 1'b0;
		Yinport_19_ <= 1'b0;
		Yinport_20_ <= 1'b0;
		Yinport_21_ <= 1'b0;
		Yinport_22_ <= 1'b0;
		Yinport_23_ <= 1'b0;
		Yinport_24_ <= 1'b0;
		Yinport_25_ <= 1'b0;
		Yinport_26_ <= 1'b0;
		Yinport_27_ <= 1'b0;
		Yinport_28_ <= 1'b0;
		Yinport_29_ <= 1'b0;
		Yinport_30_ <= 1'b0;
		Yinport_31_ <= 1'b0;
		Uinport_0_ <= 1'b0;
		Uinport_1_ <= 1'b0;
		Uinport_2_ <= 1'b0;
		Uinport_3_ <= 1'b0;
		Uinport_4_ <= 1'b0;
		Uinport_5_ <= 1'b0;
		Uinport_6_ <= 1'b0;
		Uinport_7_ <= 1'b0;
		Uinport_8_ <= 1'b0;
		Uinport_9_ <= 1'b0;
		Uinport_10_ <= 1'b0;
		Uinport_11_ <= 1'b0;
		Uinport_12_ <= 1'b0;
		Uinport_13_ <= 1'b0;
		Uinport_14_ <= 1'b0;
		Uinport_15_ <= 1'b0;
		Uinport_16_ <= 1'b0;
		Uinport_17_ <= 1'b0;
		Uinport_18_ <= 1'b0;
		Uinport_19_ <= 1'b0;
		Uinport_20_ <= 1'b0;
		Uinport_21_ <= 1'b0;
		Uinport_22_ <= 1'b0;
		Uinport_23_ <= 1'b0;
		Uinport_24_ <= 1'b0;
		Uinport_25_ <= 1'b0;
		Uinport_26_ <= 1'b0;
		Uinport_27_ <= 1'b0;
		Uinport_28_ <= 1'b0;
		Uinport_29_ <= 1'b0;
		Uinport_30_ <= 1'b0;
		Uinport_31_ <= 1'b0;
		Aport_0_ <= 1'b0;
		Aport_1_ <= 1'b0;
		Aport_2_ <= 1'b0;
		Aport_3_ <= 1'b0;
		Aport_4_ <= 1'b0;
		Aport_5_ <= 1'b0;
		Aport_6_ <= 1'b0;
		Aport_7_ <= 1'b0;
		Aport_8_ <= 1'b0;
		Aport_9_ <= 1'b0;
		Aport_10_ <= 1'b0;
		Aport_11_ <= 1'b0;
		Aport_12_ <= 1'b0;
		Aport_13_ <= 1'b0;
		Aport_14_ <= 1'b0;
		Aport_15_ <= 1'b0;
		Aport_16_ <= 1'b0;
		Aport_17_ <= 1'b0;
		Aport_18_ <= 1'b0;
		Aport_19_ <= 1'b0;
		Aport_20_ <= 1'b0;
		Aport_21_ <= 1'b0;
		Aport_22_ <= 1'b0;
		Aport_23_ <= 1'b0;
		Aport_24_ <= 1'b0;
		Aport_25_ <= 1'b0;
		Aport_26_ <= 1'b0;
		Aport_27_ <= 1'b0;
		Aport_28_ <= 1'b0;
		Aport_29_ <= 1'b0;
		Aport_30_ <= 1'b0;
		Aport_31_ <= 1'b0;
		DXport_0_ <= 1'b0;
		DXport_1_ <= 1'b0;
		DXport_2_ <= 1'b0;
		DXport_3_ <= 1'b0;
		DXport_4_ <= 1'b0;
		DXport_5_ <= 1'b0;
		DXport_6_ <= 1'b0;
		DXport_7_ <= 1'b0;
		DXport_8_ <= 1'b0;
		DXport_9_ <= 1'b0;
		DXport_10_ <= 1'b0;
		DXport_11_ <= 1'b0;
		DXport_12_ <= 1'b0;
		DXport_13_ <= 1'b0;
		DXport_14_ <= 1'b0;
		DXport_15_ <= 1'b0;
		DXport_16_ <= 1'b0;
		DXport_17_ <= 1'b0;
		DXport_18_ <= 1'b0;
		DXport_19_ <= 1'b0;
		DXport_20_ <= 1'b0;
		DXport_21_ <= 1'b0;
		DXport_22_ <= 1'b0;
		DXport_23_ <= 1'b0;
		DXport_24_ <= 1'b0;
		DXport_25_ <= 1'b0;
		DXport_26_ <= 1'b0;
		DXport_27_ <= 1'b0;
		DXport_28_ <= 1'b0;
		DXport_29_ <= 1'b0;
		DXport_30_ <= 1'b0;
		DXport_31_ <= 1'b0;
		reset <= 1'b0;

		Xoutport_0__flag[0] <= 1'b0;
		Xoutport_1__flag[0] <= 1'b0;
		Xoutport_2__flag[0] <= 1'b0;
		Xoutport_3__flag[0] <= 1'b0;
		Xoutport_4__flag[0] <= 1'b0;
		Xoutport_5__flag[0] <= 1'b0;
		Xoutport_6__flag[0] <= 1'b0;
		Xoutport_7__flag[0] <= 1'b0;
		Xoutport_8__flag[0] <= 1'b0;
		Xoutport_9__flag[0] <= 1'b0;
		Xoutport_10__flag[0] <= 1'b0;
		Xoutport_11__flag[0] <= 1'b0;
		Xoutport_12__flag[0] <= 1'b0;
		Xoutport_13__flag[0] <= 1'b0;
		Xoutport_14__flag[0] <= 1'b0;
		Xoutport_15__flag[0] <= 1'b0;
		Xoutport_16__flag[0] <= 1'b0;
		Xoutport_17__flag[0] <= 1'b0;
		Xoutport_18__flag[0] <= 1'b0;
		Xoutport_19__flag[0] <= 1'b0;
		Xoutport_20__flag[0] <= 1'b0;
		Xoutport_21__flag[0] <= 1'b0;
		Xoutport_22__flag[0] <= 1'b0;
		Xoutport_23__flag[0] <= 1'b0;
		Xoutport_24__flag[0] <= 1'b0;
		Xoutport_25__flag[0] <= 1'b0;
		Xoutport_26__flag[0] <= 1'b0;
		Xoutport_27__flag[0] <= 1'b0;
		Xoutport_28__flag[0] <= 1'b0;
		Xoutport_29__flag[0] <= 1'b0;
		Xoutport_30__flag[0] <= 1'b0;
		Xoutport_31__flag[0] <= 1'b0;
		Youtport_0__flag[0] <= 1'b0;
		Youtport_1__flag[0] <= 1'b0;
		Youtport_2__flag[0] <= 1'b0;
		Youtport_3__flag[0] <= 1'b0;
		Youtport_4__flag[0] <= 1'b0;
		Youtport_5__flag[0] <= 1'b0;
		Youtport_6__flag[0] <= 1'b0;
		Youtport_7__flag[0] <= 1'b0;
		Youtport_8__flag[0] <= 1'b0;
		Youtport_9__flag[0] <= 1'b0;
		Youtport_10__flag[0] <= 1'b0;
		Youtport_11__flag[0] <= 1'b0;
		Youtport_12__flag[0] <= 1'b0;
		Youtport_13__flag[0] <= 1'b0;
		Youtport_14__flag[0] <= 1'b0;
		Youtport_15__flag[0] <= 1'b0;
		Youtport_16__flag[0] <= 1'b0;
		Youtport_17__flag[0] <= 1'b0;
		Youtport_18__flag[0] <= 1'b0;
		Youtport_19__flag[0] <= 1'b0;
		Youtport_20__flag[0] <= 1'b0;
		Youtport_21__flag[0] <= 1'b0;
		Youtport_22__flag[0] <= 1'b0;
		Youtport_23__flag[0] <= 1'b0;
		Youtport_24__flag[0] <= 1'b0;
		Youtport_25__flag[0] <= 1'b0;
		Youtport_26__flag[0] <= 1'b0;
		Youtport_27__flag[0] <= 1'b0;
		Youtport_28__flag[0] <= 1'b0;
		Youtport_29__flag[0] <= 1'b0;
		Youtport_30__flag[0] <= 1'b0;
		Youtport_31__flag[0] <= 1'b0;
		Uoutport_0__flag[0] <= 1'b0;
		Uoutport_1__flag[0] <= 1'b0;
		Uoutport_2__flag[0] <= 1'b0;
		Uoutport_3__flag[0] <= 1'b0;
		Uoutport_4__flag[0] <= 1'b0;
		Uoutport_5__flag[0] <= 1'b0;
		Uoutport_6__flag[0] <= 1'b0;
		Uoutport_7__flag[0] <= 1'b0;
		Uoutport_8__flag[0] <= 1'b0;
		Uoutport_9__flag[0] <= 1'b0;
		Uoutport_10__flag[0] <= 1'b0;
		Uoutport_11__flag[0] <= 1'b0;
		Uoutport_12__flag[0] <= 1'b0;
		Uoutport_13__flag[0] <= 1'b0;
		Uoutport_14__flag[0] <= 1'b0;
		Uoutport_15__flag[0] <= 1'b0;
		Uoutport_16__flag[0] <= 1'b0;
		Uoutport_17__flag[0] <= 1'b0;
		Uoutport_18__flag[0] <= 1'b0;
		Uoutport_19__flag[0] <= 1'b0;
		Uoutport_20__flag[0] <= 1'b0;
		Uoutport_21__flag[0] <= 1'b0;
		Uoutport_22__flag[0] <= 1'b0;
		Uoutport_23__flag[0] <= 1'b0;
		Uoutport_24__flag[0] <= 1'b0;
		Uoutport_25__flag[0] <= 1'b0;
		Uoutport_26__flag[0] <= 1'b0;
		Uoutport_27__flag[0] <= 1'b0;
		Uoutport_28__flag[0] <= 1'b0;
		Uoutport_29__flag[0] <= 1'b0;
		Uoutport_30__flag[0] <= 1'b0;
		Uoutport_31__flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge clk[0]) begin
		Xinport_0_ <= $random;
		Xinport_1_ <= $random;
		Xinport_2_ <= $random;
		Xinport_3_ <= $random;
		Xinport_4_ <= $random;
		Xinport_5_ <= $random;
		Xinport_6_ <= $random;
		Xinport_7_ <= $random;
		Xinport_8_ <= $random;
		Xinport_9_ <= $random;
		Xinport_10_ <= $random;
		Xinport_11_ <= $random;
		Xinport_12_ <= $random;
		Xinport_13_ <= $random;
		Xinport_14_ <= $random;
		Xinport_15_ <= $random;
		Xinport_16_ <= $random;
		Xinport_17_ <= $random;
		Xinport_18_ <= $random;
		Xinport_19_ <= $random;
		Xinport_20_ <= $random;
		Xinport_21_ <= $random;
		Xinport_22_ <= $random;
		Xinport_23_ <= $random;
		Xinport_24_ <= $random;
		Xinport_25_ <= $random;
		Xinport_26_ <= $random;
		Xinport_27_ <= $random;
		Xinport_28_ <= $random;
		Xinport_29_ <= $random;
		Xinport_30_ <= $random;
		Xinport_31_ <= $random;
		Yinport_0_ <= $random;
		Yinport_1_ <= $random;
		Yinport_2_ <= $random;
		Yinport_3_ <= $random;
		Yinport_4_ <= $random;
		Yinport_5_ <= $random;
		Yinport_6_ <= $random;
		Yinport_7_ <= $random;
		Yinport_8_ <= $random;
		Yinport_9_ <= $random;
		Yinport_10_ <= $random;
		Yinport_11_ <= $random;
		Yinport_12_ <= $random;
		Yinport_13_ <= $random;
		Yinport_14_ <= $random;
		Yinport_15_ <= $random;
		Yinport_16_ <= $random;
		Yinport_17_ <= $random;
		Yinport_18_ <= $random;
		Yinport_19_ <= $random;
		Yinport_20_ <= $random;
		Yinport_21_ <= $random;
		Yinport_22_ <= $random;
		Yinport_23_ <= $random;
		Yinport_24_ <= $random;
		Yinport_25_ <= $random;
		Yinport_26_ <= $random;
		Yinport_27_ <= $random;
		Yinport_28_ <= $random;
		Yinport_29_ <= $random;
		Yinport_30_ <= $random;
		Yinport_31_ <= $random;
		Uinport_0_ <= $random;
		Uinport_1_ <= $random;
		Uinport_2_ <= $random;
		Uinport_3_ <= $random;
		Uinport_4_ <= $random;
		Uinport_5_ <= $random;
		Uinport_6_ <= $random;
		Uinport_7_ <= $random;
		Uinport_8_ <= $random;
		Uinport_9_ <= $random;
		Uinport_10_ <= $random;
		Uinport_11_ <= $random;
		Uinport_12_ <= $random;
		Uinport_13_ <= $random;
		Uinport_14_ <= $random;
		Uinport_15_ <= $random;
		Uinport_16_ <= $random;
		Uinport_17_ <= $random;
		Uinport_18_ <= $random;
		Uinport_19_ <= $random;
		Uinport_20_ <= $random;
		Uinport_21_ <= $random;
		Uinport_22_ <= $random;
		Uinport_23_ <= $random;
		Uinport_24_ <= $random;
		Uinport_25_ <= $random;
		Uinport_26_ <= $random;
		Uinport_27_ <= $random;
		Uinport_28_ <= $random;
		Uinport_29_ <= $random;
		Uinport_30_ <= $random;
		Uinport_31_ <= $random;
		Aport_0_ <= $random;
		Aport_1_ <= $random;
		Aport_2_ <= $random;
		Aport_3_ <= $random;
		Aport_4_ <= $random;
		Aport_5_ <= $random;
		Aport_6_ <= $random;
		Aport_7_ <= $random;
		Aport_8_ <= $random;
		Aport_9_ <= $random;
		Aport_10_ <= $random;
		Aport_11_ <= $random;
		Aport_12_ <= $random;
		Aport_13_ <= $random;
		Aport_14_ <= $random;
		Aport_15_ <= $random;
		Aport_16_ <= $random;
		Aport_17_ <= $random;
		Aport_18_ <= $random;
		Aport_19_ <= $random;
		Aport_20_ <= $random;
		Aport_21_ <= $random;
		Aport_22_ <= $random;
		Aport_23_ <= $random;
		Aport_24_ <= $random;
		Aport_25_ <= $random;
		Aport_26_ <= $random;
		Aport_27_ <= $random;
		Aport_28_ <= $random;
		Aport_29_ <= $random;
		Aport_30_ <= $random;
		Aport_31_ <= $random;
		DXport_0_ <= $random;
		DXport_1_ <= $random;
		DXport_2_ <= $random;
		DXport_3_ <= $random;
		DXport_4_ <= $random;
		DXport_5_ <= $random;
		DXport_6_ <= $random;
		DXport_7_ <= $random;
		DXport_8_ <= $random;
		DXport_9_ <= $random;
		DXport_10_ <= $random;
		DXport_11_ <= $random;
		DXport_12_ <= $random;
		DXport_13_ <= $random;
		DXport_14_ <= $random;
		DXport_15_ <= $random;
		DXport_16_ <= $random;
		DXport_17_ <= $random;
		DXport_18_ <= $random;
		DXport_19_ <= $random;
		DXport_20_ <= $random;
		DXport_21_ <= $random;
		DXport_22_ <= $random;
		DXport_23_ <= $random;
		DXport_24_ <= $random;
		DXport_25_ <= $random;
		DXport_26_ <= $random;
		DXport_27_ <= $random;
		DXport_28_ <= $random;
		DXport_29_ <= $random;
		DXport_30_ <= $random;
		DXport_31_ <= $random;
		reset <= $random;
	end

// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge clk[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else 
begin
			if(!(Xoutport_0__gfpga === Xoutport_0__bench) && !(Xoutport_0__bench === 1'bx)) begin
				Xoutport_0__flag <= 1'b1;
			end else begin
				Xoutport_0__flag<= 1'b0;
			end
			if(!(Xoutport_1__gfpga === Xoutport_1__bench) && !(Xoutport_1__bench === 1'bx)) begin
				Xoutport_1__flag <= 1'b1;
			end else begin
				Xoutport_1__flag<= 1'b0;
			end
			if(!(Xoutport_2__gfpga === Xoutport_2__bench) && !(Xoutport_2__bench === 1'bx)) begin
				Xoutport_2__flag <= 1'b1;
			end else begin
				Xoutport_2__flag<= 1'b0;
			end
			if(!(Xoutport_3__gfpga === Xoutport_3__bench) && !(Xoutport_3__bench === 1'bx)) begin
				Xoutport_3__flag <= 1'b1;
			end else begin
				Xoutport_3__flag<= 1'b0;
			end
			if(!(Xoutport_4__gfpga === Xoutport_4__bench) && !(Xoutport_4__bench === 1'bx)) begin
				Xoutport_4__flag <= 1'b1;
			end else begin
				Xoutport_4__flag<= 1'b0;
			end
			if(!(Xoutport_5__gfpga === Xoutport_5__bench) && !(Xoutport_5__bench === 1'bx)) begin
				Xoutport_5__flag <= 1'b1;
			end else begin
				Xoutport_5__flag<= 1'b0;
			end
			if(!(Xoutport_6__gfpga === Xoutport_6__bench) && !(Xoutport_6__bench === 1'bx)) begin
				Xoutport_6__flag <= 1'b1;
			end else begin
				Xoutport_6__flag<= 1'b0;
			end
			if(!(Xoutport_7__gfpga === Xoutport_7__bench) && !(Xoutport_7__bench === 1'bx)) begin
				Xoutport_7__flag <= 1'b1;
			end else begin
				Xoutport_7__flag<= 1'b0;
			end
			if(!(Xoutport_8__gfpga === Xoutport_8__bench) && !(Xoutport_8__bench === 1'bx)) begin
				Xoutport_8__flag <= 1'b1;
			end else begin
				Xoutport_8__flag<= 1'b0;
			end
			if(!(Xoutport_9__gfpga === Xoutport_9__bench) && !(Xoutport_9__bench === 1'bx)) begin
				Xoutport_9__flag <= 1'b1;
			end else begin
				Xoutport_9__flag<= 1'b0;
			end
			if(!(Xoutport_10__gfpga === Xoutport_10__bench) && !(Xoutport_10__bench === 1'bx)) begin
				Xoutport_10__flag <= 1'b1;
			end else begin
				Xoutport_10__flag<= 1'b0;
			end
			if(!(Xoutport_11__gfpga === Xoutport_11__bench) && !(Xoutport_11__bench === 1'bx)) begin
				Xoutport_11__flag <= 1'b1;
			end else begin
				Xoutport_11__flag<= 1'b0;
			end
			if(!(Xoutport_12__gfpga === Xoutport_12__bench) && !(Xoutport_12__bench === 1'bx)) begin
				Xoutport_12__flag <= 1'b1;
			end else begin
				Xoutport_12__flag<= 1'b0;
			end
			if(!(Xoutport_13__gfpga === Xoutport_13__bench) && !(Xoutport_13__bench === 1'bx)) begin
				Xoutport_13__flag <= 1'b1;
			end else begin
				Xoutport_13__flag<= 1'b0;
			end
			if(!(Xoutport_14__gfpga === Xoutport_14__bench) && !(Xoutport_14__bench === 1'bx)) begin
				Xoutport_14__flag <= 1'b1;
			end else begin
				Xoutport_14__flag<= 1'b0;
			end
			if(!(Xoutport_15__gfpga === Xoutport_15__bench) && !(Xoutport_15__bench === 1'bx)) begin
				Xoutport_15__flag <= 1'b1;
			end else begin
				Xoutport_15__flag<= 1'b0;
			end
			if(!(Xoutport_16__gfpga === Xoutport_16__bench) && !(Xoutport_16__bench === 1'bx)) begin
				Xoutport_16__flag <= 1'b1;
			end else begin
				Xoutport_16__flag<= 1'b0;
			end
			if(!(Xoutport_17__gfpga === Xoutport_17__bench) && !(Xoutport_17__bench === 1'bx)) begin
				Xoutport_17__flag <= 1'b1;
			end else begin
				Xoutport_17__flag<= 1'b0;
			end
			if(!(Xoutport_18__gfpga === Xoutport_18__bench) && !(Xoutport_18__bench === 1'bx)) begin
				Xoutport_18__flag <= 1'b1;
			end else begin
				Xoutport_18__flag<= 1'b0;
			end
			if(!(Xoutport_19__gfpga === Xoutport_19__bench) && !(Xoutport_19__bench === 1'bx)) begin
				Xoutport_19__flag <= 1'b1;
			end else begin
				Xoutport_19__flag<= 1'b0;
			end
			if(!(Xoutport_20__gfpga === Xoutport_20__bench) && !(Xoutport_20__bench === 1'bx)) begin
				Xoutport_20__flag <= 1'b1;
			end else begin
				Xoutport_20__flag<= 1'b0;
			end
			if(!(Xoutport_21__gfpga === Xoutport_21__bench) && !(Xoutport_21__bench === 1'bx)) begin
				Xoutport_21__flag <= 1'b1;
			end else begin
				Xoutport_21__flag<= 1'b0;
			end
			if(!(Xoutport_22__gfpga === Xoutport_22__bench) && !(Xoutport_22__bench === 1'bx)) begin
				Xoutport_22__flag <= 1'b1;
			end else begin
				Xoutport_22__flag<= 1'b0;
			end
			if(!(Xoutport_23__gfpga === Xoutport_23__bench) && !(Xoutport_23__bench === 1'bx)) begin
				Xoutport_23__flag <= 1'b1;
			end else begin
				Xoutport_23__flag<= 1'b0;
			end
			if(!(Xoutport_24__gfpga === Xoutport_24__bench) && !(Xoutport_24__bench === 1'bx)) begin
				Xoutport_24__flag <= 1'b1;
			end else begin
				Xoutport_24__flag<= 1'b0;
			end
			if(!(Xoutport_25__gfpga === Xoutport_25__bench) && !(Xoutport_25__bench === 1'bx)) begin
				Xoutport_25__flag <= 1'b1;
			end else begin
				Xoutport_25__flag<= 1'b0;
			end
			if(!(Xoutport_26__gfpga === Xoutport_26__bench) && !(Xoutport_26__bench === 1'bx)) begin
				Xoutport_26__flag <= 1'b1;
			end else begin
				Xoutport_26__flag<= 1'b0;
			end
			if(!(Xoutport_27__gfpga === Xoutport_27__bench) && !(Xoutport_27__bench === 1'bx)) begin
				Xoutport_27__flag <= 1'b1;
			end else begin
				Xoutport_27__flag<= 1'b0;
			end
			if(!(Xoutport_28__gfpga === Xoutport_28__bench) && !(Xoutport_28__bench === 1'bx)) begin
				Xoutport_28__flag <= 1'b1;
			end else begin
				Xoutport_28__flag<= 1'b0;
			end
			if(!(Xoutport_29__gfpga === Xoutport_29__bench) && !(Xoutport_29__bench === 1'bx)) begin
				Xoutport_29__flag <= 1'b1;
			end else begin
				Xoutport_29__flag<= 1'b0;
			end
			if(!(Xoutport_30__gfpga === Xoutport_30__bench) && !(Xoutport_30__bench === 1'bx)) begin
				Xoutport_30__flag <= 1'b1;
			end else begin
				Xoutport_30__flag<= 1'b0;
			end
			if(!(Xoutport_31__gfpga === Xoutport_31__bench) && !(Xoutport_31__bench === 1'bx)) begin
				Xoutport_31__flag <= 1'b1;
			end else begin
				Xoutport_31__flag<= 1'b0;
			end
			if(!(Youtport_0__gfpga === Youtport_0__bench) && !(Youtport_0__bench === 1'bx)) begin
				Youtport_0__flag <= 1'b1;
			end else begin
				Youtport_0__flag<= 1'b0;
			end
			if(!(Youtport_1__gfpga === Youtport_1__bench) && !(Youtport_1__bench === 1'bx)) begin
				Youtport_1__flag <= 1'b1;
			end else begin
				Youtport_1__flag<= 1'b0;
			end
			if(!(Youtport_2__gfpga === Youtport_2__bench) && !(Youtport_2__bench === 1'bx)) begin
				Youtport_2__flag <= 1'b1;
			end else begin
				Youtport_2__flag<= 1'b0;
			end
			if(!(Youtport_3__gfpga === Youtport_3__bench) && !(Youtport_3__bench === 1'bx)) begin
				Youtport_3__flag <= 1'b1;
			end else begin
				Youtport_3__flag<= 1'b0;
			end
			if(!(Youtport_4__gfpga === Youtport_4__bench) && !(Youtport_4__bench === 1'bx)) begin
				Youtport_4__flag <= 1'b1;
			end else begin
				Youtport_4__flag<= 1'b0;
			end
			if(!(Youtport_5__gfpga === Youtport_5__bench) && !(Youtport_5__bench === 1'bx)) begin
				Youtport_5__flag <= 1'b1;
			end else begin
				Youtport_5__flag<= 1'b0;
			end
			if(!(Youtport_6__gfpga === Youtport_6__bench) && !(Youtport_6__bench === 1'bx)) begin
				Youtport_6__flag <= 1'b1;
			end else begin
				Youtport_6__flag<= 1'b0;
			end
			if(!(Youtport_7__gfpga === Youtport_7__bench) && !(Youtport_7__bench === 1'bx)) begin
				Youtport_7__flag <= 1'b1;
			end else begin
				Youtport_7__flag<= 1'b0;
			end
			if(!(Youtport_8__gfpga === Youtport_8__bench) && !(Youtport_8__bench === 1'bx)) begin
				Youtport_8__flag <= 1'b1;
			end else begin
				Youtport_8__flag<= 1'b0;
			end
			if(!(Youtport_9__gfpga === Youtport_9__bench) && !(Youtport_9__bench === 1'bx)) begin
				Youtport_9__flag <= 1'b1;
			end else begin
				Youtport_9__flag<= 1'b0;
			end
			if(!(Youtport_10__gfpga === Youtport_10__bench) && !(Youtport_10__bench === 1'bx)) begin
				Youtport_10__flag <= 1'b1;
			end else begin
				Youtport_10__flag<= 1'b0;
			end
			if(!(Youtport_11__gfpga === Youtport_11__bench) && !(Youtport_11__bench === 1'bx)) begin
				Youtport_11__flag <= 1'b1;
			end else begin
				Youtport_11__flag<= 1'b0;
			end
			if(!(Youtport_12__gfpga === Youtport_12__bench) && !(Youtport_12__bench === 1'bx)) begin
				Youtport_12__flag <= 1'b1;
			end else begin
				Youtport_12__flag<= 1'b0;
			end
			if(!(Youtport_13__gfpga === Youtport_13__bench) && !(Youtport_13__bench === 1'bx)) begin
				Youtport_13__flag <= 1'b1;
			end else begin
				Youtport_13__flag<= 1'b0;
			end
			if(!(Youtport_14__gfpga === Youtport_14__bench) && !(Youtport_14__bench === 1'bx)) begin
				Youtport_14__flag <= 1'b1;
			end else begin
				Youtport_14__flag<= 1'b0;
			end
			if(!(Youtport_15__gfpga === Youtport_15__bench) && !(Youtport_15__bench === 1'bx)) begin
				Youtport_15__flag <= 1'b1;
			end else begin
				Youtport_15__flag<= 1'b0;
			end
			if(!(Youtport_16__gfpga === Youtport_16__bench) && !(Youtport_16__bench === 1'bx)) begin
				Youtport_16__flag <= 1'b1;
			end else begin
				Youtport_16__flag<= 1'b0;
			end
			if(!(Youtport_17__gfpga === Youtport_17__bench) && !(Youtport_17__bench === 1'bx)) begin
				Youtport_17__flag <= 1'b1;
			end else begin
				Youtport_17__flag<= 1'b0;
			end
			if(!(Youtport_18__gfpga === Youtport_18__bench) && !(Youtport_18__bench === 1'bx)) begin
				Youtport_18__flag <= 1'b1;
			end else begin
				Youtport_18__flag<= 1'b0;
			end
			if(!(Youtport_19__gfpga === Youtport_19__bench) && !(Youtport_19__bench === 1'bx)) begin
				Youtport_19__flag <= 1'b1;
			end else begin
				Youtport_19__flag<= 1'b0;
			end
			if(!(Youtport_20__gfpga === Youtport_20__bench) && !(Youtport_20__bench === 1'bx)) begin
				Youtport_20__flag <= 1'b1;
			end else begin
				Youtport_20__flag<= 1'b0;
			end
			if(!(Youtport_21__gfpga === Youtport_21__bench) && !(Youtport_21__bench === 1'bx)) begin
				Youtport_21__flag <= 1'b1;
			end else begin
				Youtport_21__flag<= 1'b0;
			end
			if(!(Youtport_22__gfpga === Youtport_22__bench) && !(Youtport_22__bench === 1'bx)) begin
				Youtport_22__flag <= 1'b1;
			end else begin
				Youtport_22__flag<= 1'b0;
			end
			if(!(Youtport_23__gfpga === Youtport_23__bench) && !(Youtport_23__bench === 1'bx)) begin
				Youtport_23__flag <= 1'b1;
			end else begin
				Youtport_23__flag<= 1'b0;
			end
			if(!(Youtport_24__gfpga === Youtport_24__bench) && !(Youtport_24__bench === 1'bx)) begin
				Youtport_24__flag <= 1'b1;
			end else begin
				Youtport_24__flag<= 1'b0;
			end
			if(!(Youtport_25__gfpga === Youtport_25__bench) && !(Youtport_25__bench === 1'bx)) begin
				Youtport_25__flag <= 1'b1;
			end else begin
				Youtport_25__flag<= 1'b0;
			end
			if(!(Youtport_26__gfpga === Youtport_26__bench) && !(Youtport_26__bench === 1'bx)) begin
				Youtport_26__flag <= 1'b1;
			end else begin
				Youtport_26__flag<= 1'b0;
			end
			if(!(Youtport_27__gfpga === Youtport_27__bench) && !(Youtport_27__bench === 1'bx)) begin
				Youtport_27__flag <= 1'b1;
			end else begin
				Youtport_27__flag<= 1'b0;
			end
			if(!(Youtport_28__gfpga === Youtport_28__bench) && !(Youtport_28__bench === 1'bx)) begin
				Youtport_28__flag <= 1'b1;
			end else begin
				Youtport_28__flag<= 1'b0;
			end
			if(!(Youtport_29__gfpga === Youtport_29__bench) && !(Youtport_29__bench === 1'bx)) begin
				Youtport_29__flag <= 1'b1;
			end else begin
				Youtport_29__flag<= 1'b0;
			end
			if(!(Youtport_30__gfpga === Youtport_30__bench) && !(Youtport_30__bench === 1'bx)) begin
				Youtport_30__flag <= 1'b1;
			end else begin
				Youtport_30__flag<= 1'b0;
			end
			if(!(Youtport_31__gfpga === Youtport_31__bench) && !(Youtport_31__bench === 1'bx)) begin
				Youtport_31__flag <= 1'b1;
			end else begin
				Youtport_31__flag<= 1'b0;
			end
			if(!(Uoutport_0__gfpga === Uoutport_0__bench) && !(Uoutport_0__bench === 1'bx)) begin
				Uoutport_0__flag <= 1'b1;
			end else begin
				Uoutport_0__flag<= 1'b0;
			end
			if(!(Uoutport_1__gfpga === Uoutport_1__bench) && !(Uoutport_1__bench === 1'bx)) begin
				Uoutport_1__flag <= 1'b1;
			end else begin
				Uoutport_1__flag<= 1'b0;
			end
			if(!(Uoutport_2__gfpga === Uoutport_2__bench) && !(Uoutport_2__bench === 1'bx)) begin
				Uoutport_2__flag <= 1'b1;
			end else begin
				Uoutport_2__flag<= 1'b0;
			end
			if(!(Uoutport_3__gfpga === Uoutport_3__bench) && !(Uoutport_3__bench === 1'bx)) begin
				Uoutport_3__flag <= 1'b1;
			end else begin
				Uoutport_3__flag<= 1'b0;
			end
			if(!(Uoutport_4__gfpga === Uoutport_4__bench) && !(Uoutport_4__bench === 1'bx)) begin
				Uoutport_4__flag <= 1'b1;
			end else begin
				Uoutport_4__flag<= 1'b0;
			end
			if(!(Uoutport_5__gfpga === Uoutport_5__bench) && !(Uoutport_5__bench === 1'bx)) begin
				Uoutport_5__flag <= 1'b1;
			end else begin
				Uoutport_5__flag<= 1'b0;
			end
			if(!(Uoutport_6__gfpga === Uoutport_6__bench) && !(Uoutport_6__bench === 1'bx)) begin
				Uoutport_6__flag <= 1'b1;
			end else begin
				Uoutport_6__flag<= 1'b0;
			end
			if(!(Uoutport_7__gfpga === Uoutport_7__bench) && !(Uoutport_7__bench === 1'bx)) begin
				Uoutport_7__flag <= 1'b1;
			end else begin
				Uoutport_7__flag<= 1'b0;
			end
			if(!(Uoutport_8__gfpga === Uoutport_8__bench) && !(Uoutport_8__bench === 1'bx)) begin
				Uoutport_8__flag <= 1'b1;
			end else begin
				Uoutport_8__flag<= 1'b0;
			end
			if(!(Uoutport_9__gfpga === Uoutport_9__bench) && !(Uoutport_9__bench === 1'bx)) begin
				Uoutport_9__flag <= 1'b1;
			end else begin
				Uoutport_9__flag<= 1'b0;
			end
			if(!(Uoutport_10__gfpga === Uoutport_10__bench) && !(Uoutport_10__bench === 1'bx)) begin
				Uoutport_10__flag <= 1'b1;
			end else begin
				Uoutport_10__flag<= 1'b0;
			end
			if(!(Uoutport_11__gfpga === Uoutport_11__bench) && !(Uoutport_11__bench === 1'bx)) begin
				Uoutport_11__flag <= 1'b1;
			end else begin
				Uoutport_11__flag<= 1'b0;
			end
			if(!(Uoutport_12__gfpga === Uoutport_12__bench) && !(Uoutport_12__bench === 1'bx)) begin
				Uoutport_12__flag <= 1'b1;
			end else begin
				Uoutport_12__flag<= 1'b0;
			end
			if(!(Uoutport_13__gfpga === Uoutport_13__bench) && !(Uoutport_13__bench === 1'bx)) begin
				Uoutport_13__flag <= 1'b1;
			end else begin
				Uoutport_13__flag<= 1'b0;
			end
			if(!(Uoutport_14__gfpga === Uoutport_14__bench) && !(Uoutport_14__bench === 1'bx)) begin
				Uoutport_14__flag <= 1'b1;
			end else begin
				Uoutport_14__flag<= 1'b0;
			end
			if(!(Uoutport_15__gfpga === Uoutport_15__bench) && !(Uoutport_15__bench === 1'bx)) begin
				Uoutport_15__flag <= 1'b1;
			end else begin
				Uoutport_15__flag<= 1'b0;
			end
			if(!(Uoutport_16__gfpga === Uoutport_16__bench) && !(Uoutport_16__bench === 1'bx)) begin
				Uoutport_16__flag <= 1'b1;
			end else begin
				Uoutport_16__flag<= 1'b0;
			end
			if(!(Uoutport_17__gfpga === Uoutport_17__bench) && !(Uoutport_17__bench === 1'bx)) begin
				Uoutport_17__flag <= 1'b1;
			end else begin
				Uoutport_17__flag<= 1'b0;
			end
			if(!(Uoutport_18__gfpga === Uoutport_18__bench) && !(Uoutport_18__bench === 1'bx)) begin
				Uoutport_18__flag <= 1'b1;
			end else begin
				Uoutport_18__flag<= 1'b0;
			end
			if(!(Uoutport_19__gfpga === Uoutport_19__bench) && !(Uoutport_19__bench === 1'bx)) begin
				Uoutport_19__flag <= 1'b1;
			end else begin
				Uoutport_19__flag<= 1'b0;
			end
			if(!(Uoutport_20__gfpga === Uoutport_20__bench) && !(Uoutport_20__bench === 1'bx)) begin
				Uoutport_20__flag <= 1'b1;
			end else begin
				Uoutport_20__flag<= 1'b0;
			end
			if(!(Uoutport_21__gfpga === Uoutport_21__bench) && !(Uoutport_21__bench === 1'bx)) begin
				Uoutport_21__flag <= 1'b1;
			end else begin
				Uoutport_21__flag<= 1'b0;
			end
			if(!(Uoutport_22__gfpga === Uoutport_22__bench) && !(Uoutport_22__bench === 1'bx)) begin
				Uoutport_22__flag <= 1'b1;
			end else begin
				Uoutport_22__flag<= 1'b0;
			end
			if(!(Uoutport_23__gfpga === Uoutport_23__bench) && !(Uoutport_23__bench === 1'bx)) begin
				Uoutport_23__flag <= 1'b1;
			end else begin
				Uoutport_23__flag<= 1'b0;
			end
			if(!(Uoutport_24__gfpga === Uoutport_24__bench) && !(Uoutport_24__bench === 1'bx)) begin
				Uoutport_24__flag <= 1'b1;
			end else begin
				Uoutport_24__flag<= 1'b0;
			end
			if(!(Uoutport_25__gfpga === Uoutport_25__bench) && !(Uoutport_25__bench === 1'bx)) begin
				Uoutport_25__flag <= 1'b1;
			end else begin
				Uoutport_25__flag<= 1'b0;
			end
			if(!(Uoutport_26__gfpga === Uoutport_26__bench) && !(Uoutport_26__bench === 1'bx)) begin
				Uoutport_26__flag <= 1'b1;
			end else begin
				Uoutport_26__flag<= 1'b0;
			end
			if(!(Uoutport_27__gfpga === Uoutport_27__bench) && !(Uoutport_27__bench === 1'bx)) begin
				Uoutport_27__flag <= 1'b1;
			end else begin
				Uoutport_27__flag<= 1'b0;
			end
			if(!(Uoutport_28__gfpga === Uoutport_28__bench) && !(Uoutport_28__bench === 1'bx)) begin
				Uoutport_28__flag <= 1'b1;
			end else begin
				Uoutport_28__flag<= 1'b0;
			end
			if(!(Uoutport_29__gfpga === Uoutport_29__bench) && !(Uoutport_29__bench === 1'bx)) begin
				Uoutport_29__flag <= 1'b1;
			end else begin
				Uoutport_29__flag<= 1'b0;
			end
			if(!(Uoutport_30__gfpga === Uoutport_30__bench) && !(Uoutport_30__bench === 1'bx)) begin
				Uoutport_30__flag <= 1'b1;
			end else begin
				Uoutport_30__flag<= 1'b0;
			end
			if(!(Uoutport_31__gfpga === Uoutport_31__bench) && !(Uoutport_31__bench === 1'bx)) begin
				Uoutport_31__flag <= 1'b1;
			end else begin
				Uoutport_31__flag<= 1'b0;
			end
		end
	end

	always@(posedge Xoutport_0__flag) begin
		if(Xoutport_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_1__flag) begin
		if(Xoutport_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_2__flag) begin
		if(Xoutport_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_3__flag) begin
		if(Xoutport_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_4__flag) begin
		if(Xoutport_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_5__flag) begin
		if(Xoutport_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_6__flag) begin
		if(Xoutport_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_7__flag) begin
		if(Xoutport_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_8__flag) begin
		if(Xoutport_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_9__flag) begin
		if(Xoutport_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_10__flag) begin
		if(Xoutport_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_11__flag) begin
		if(Xoutport_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_12__flag) begin
		if(Xoutport_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_13__flag) begin
		if(Xoutport_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_14__flag) begin
		if(Xoutport_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_15__flag) begin
		if(Xoutport_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_16__flag) begin
		if(Xoutport_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_17__flag) begin
		if(Xoutport_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_18__flag) begin
		if(Xoutport_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_19__flag) begin
		if(Xoutport_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_20__flag) begin
		if(Xoutport_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_21__flag) begin
		if(Xoutport_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_22__flag) begin
		if(Xoutport_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_23__flag) begin
		if(Xoutport_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_24__flag) begin
		if(Xoutport_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_25__flag) begin
		if(Xoutport_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_26__flag) begin
		if(Xoutport_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_27__flag) begin
		if(Xoutport_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_28__flag) begin
		if(Xoutport_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_29__flag) begin
		if(Xoutport_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_30__flag) begin
		if(Xoutport_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Xoutport_31__flag) begin
		if(Xoutport_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Xoutport_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_0__flag) begin
		if(Youtport_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_1__flag) begin
		if(Youtport_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_2__flag) begin
		if(Youtport_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_3__flag) begin
		if(Youtport_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_4__flag) begin
		if(Youtport_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_5__flag) begin
		if(Youtport_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_6__flag) begin
		if(Youtport_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_7__flag) begin
		if(Youtport_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_8__flag) begin
		if(Youtport_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_9__flag) begin
		if(Youtport_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_10__flag) begin
		if(Youtport_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_11__flag) begin
		if(Youtport_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_12__flag) begin
		if(Youtport_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_13__flag) begin
		if(Youtport_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_14__flag) begin
		if(Youtport_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_15__flag) begin
		if(Youtport_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_16__flag) begin
		if(Youtport_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_17__flag) begin
		if(Youtport_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_18__flag) begin
		if(Youtport_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_19__flag) begin
		if(Youtport_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_20__flag) begin
		if(Youtport_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_21__flag) begin
		if(Youtport_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_22__flag) begin
		if(Youtport_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_23__flag) begin
		if(Youtport_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_24__flag) begin
		if(Youtport_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_25__flag) begin
		if(Youtport_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_26__flag) begin
		if(Youtport_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_27__flag) begin
		if(Youtport_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_28__flag) begin
		if(Youtport_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_29__flag) begin
		if(Youtport_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_30__flag) begin
		if(Youtport_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Youtport_31__flag) begin
		if(Youtport_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Youtport_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_0__flag) begin
		if(Uoutport_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_1__flag) begin
		if(Uoutport_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_2__flag) begin
		if(Uoutport_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_3__flag) begin
		if(Uoutport_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_4__flag) begin
		if(Uoutport_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_5__flag) begin
		if(Uoutport_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_6__flag) begin
		if(Uoutport_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_7__flag) begin
		if(Uoutport_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_8__flag) begin
		if(Uoutport_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_9__flag) begin
		if(Uoutport_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_10__flag) begin
		if(Uoutport_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_11__flag) begin
		if(Uoutport_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_12__flag) begin
		if(Uoutport_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_13__flag) begin
		if(Uoutport_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_14__flag) begin
		if(Uoutport_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_15__flag) begin
		if(Uoutport_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_16__flag) begin
		if(Uoutport_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_17__flag) begin
		if(Uoutport_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_18__flag) begin
		if(Uoutport_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_19__flag) begin
		if(Uoutport_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_20__flag) begin
		if(Uoutport_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_21__flag) begin
		if(Uoutport_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_22__flag) begin
		if(Uoutport_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_23__flag) begin
		if(Uoutport_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_24__flag) begin
		if(Uoutport_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_25__flag) begin
		if(Uoutport_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_26__flag) begin
		if(Uoutport_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_27__flag) begin
		if(Uoutport_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_28__flag) begin
		if(Uoutport_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_29__flag) begin
		if(Uoutport_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_30__flag) begin
		if(Uoutport_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge Uoutport_31__flag) begin
		if(Uoutport_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on Uoutport_31__gfpga at time = %t", $realtime);
		end
	end


// ----- Begin output waveform to VCD file-------
	initial begin
		$dumpfile("diffeq_paj_convert_formal.vcd");
		$dumpvars(1, diffeq_paj_convert_top_formal_verification_random_tb);
	end
// ----- END output waveform to VCD file -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#20
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for diffeq_paj_convert_top_formal_verification_random_tb -----

